--author :Pranav Tambe
library IEEE;
use IEEE.std_logic_1164.all;
use work.CS210.all;
entity MUX_2X1 is port(I0, I1, S0 : in std_logic; -- Inputs 
                       O0 : out std_logic); -- Output 
end MUX_2X1;  
architecture STRUCTURE of MUX_2X1 is
signal SIG_S0,SIG_S1,SIG_S2:std_logic;
begin
	U0:NOT1 port map(S0,SIG_S0);--Compliment of select line S0
  	U1:AND2 port map(I0,SIG_S0,SIG_S1); --Intermediate signal SIG_S1 by AND operation (Product) I0 and Compliment of select line S0
      U2: AND2 port map(I1,S0,SIG_S2);  --Intermediate signal SIG_S2 by  AND operation (Product) on I1 and select line S0
	U3: OR2 port map(SIG_S1,SIG_S2,O0); --Output O0 by OR operation (Sum) Intermadiate signals generated by two AND gates
end STRUCTURE;   